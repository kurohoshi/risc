library ieee

entity 
