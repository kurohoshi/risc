library ieee;
   use ieee.std_logic_1164.all;

entity mult32 is
   port(
      a, b     : in std_logic_vector(31 downto 0);
    --sign     : in std_logic;
      result   : out std_logic_vector(31 downto 0)
   );
end mult32;

architecture struct of mult32 is
   --do 32-bit multiplication

   --declare any internal signals
begin
   -- do 32-bit addition
end struct;
